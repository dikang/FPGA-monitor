`ifndef __CACHES_CFG_SVH__
`define __CACHES_CFG_SVH__

`define LLSC
`define LITTLE_ENDIAN
`define ADDR_BITS    32
`define BYTE_BITS    3
`define WORD_BITS    1
`define L2_WAYS      4
`define L2_SETS      512
`define LLC_WAYS     16
`define LLC_SETS     1024
`define DMA_NOC_WIDTH    64

`endif // __CACHES_CFG_SVH__
